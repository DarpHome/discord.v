module discord
